
`uvm_analysis_imp_decl(_ip)
`uvm_analysis_imp_decl(_op)

  
  `include "evm_interface.sv"
  `include "evm_seq_item.sv"
  `include "evm_sequence.sv"
  `include "evm_sequencer.sv"
  `include "evm_driver.sv"
  `include "evm_input_monitor.sv"
  `include "evm_output_monitor.sv"
  `include "evm_active_agent.sv"
  `include "evm_passive_agent.sv"
 // `include "evm_scb.sv"
  //`include "evm_cov.sv"
  `include "evm_env.sv"
  `include "evm_test.sv"


